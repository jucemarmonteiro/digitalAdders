// Copyright {2011} {Jucemar Monteiro - jucemar.monteiro@gmail.com}
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at

// http://www.apache.org/licenses/LICENSE-2.0

// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//-----------------------------------------------------
// Design Name : rb2_mux
// File Name   : rb2_mux.v
// Function    : recomputing block for bit 3 of sum
// Coder       : Jucemar Monteiro
//-----------------------------------------------------
module  rb2_mux (s, rs);
	parameter n = 3;
	input  [n-1:0]s;
	output  rs;

	assign rs= (s[0] & s[1]) ^ s[2];
endmodule 

