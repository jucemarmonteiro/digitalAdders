// Copyright {2011} {Jucemar Monteiro - jucemar.monteiro@gmail.com}
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at

// http://www.apache.org/licenses/LICENSE-2.0

// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//
//-----------------------------------------------------
// Design Name : prop_signal
// File Name   : prop_signal.v
// Function    : Carry Propagate for 4 bit int the CLA Block
// Coder       : Jucemar Monteiro
//-----------------------------------------------------

module prop_signal (p,prop);
	parameter n=4;
	input   [n-1:0]p;
	output   prop;
	assign prop = p[0] & p[1] & p[2] & p[3];
endmodule
